module Baud_Counter #(
  parameter TIMER_BITS=10
)(
  input  wire       clk , arst_n , count_en, count_rst,
  input  wire [9:0] Load_Value,
  output wire [3:0] count 
);
  //Connection Wire
  wire done;

  //In this module, we use a timer that ticka after 1/16 of bit period specified by the baud rate
  //And another counter that counts from 0 to 15 to indicate a bit time
  //The counter output is connected to the FSM Controller inside the Tx or the Rx to take dicision upon
  //timer instantiation
  timer #(.TIMER_BITS(TIMER_BITS)) timer_inst (
    .clk(clk),
    .rst_n(arst_n),
    .rst(count_rst),
    .enable(count_en),
    .Load_Value(Load_Value),
    .done(done)
  );
  
  //Mod-16 counter instantiation
  counter counter_inst (
    .clk(clk),
    .enab(done),
    .rst_n(arst_n),
    .rst(count_rst),
    .cnt_out(count)
  );
endmodule